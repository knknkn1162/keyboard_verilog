`include "testbench.v"
`include "kb_sampling_en.v"

module kb_sampling_en_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule

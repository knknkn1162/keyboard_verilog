`include "testbench.v"
`include "shift_key.v"

module shift_key_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule

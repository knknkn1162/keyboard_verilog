`include "testbench.v"
`include "scancode2ascii.v"

module scancode2ascii_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule

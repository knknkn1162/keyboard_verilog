`include "testbench.v"
`include "recv.v"

module recv_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule

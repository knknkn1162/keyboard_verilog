`include "testbench.v"
`include "keydown.v"

module keydown_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule

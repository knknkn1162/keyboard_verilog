`include "testbench.v"
`include "keyboard.v"

module keyboard_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule

`include "testbench.v"
`include "keyboard_negedge_detector.v"

module keyboard_negedge_detector_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
